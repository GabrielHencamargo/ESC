module gnot(input a, output y);
    assign y = ~a;
endmodule